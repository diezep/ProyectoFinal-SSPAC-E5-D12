module SHIFTLEFT(
    input[31:0] OP,
    output[31:0] OPS
);

//TODO: Lógica

endmodule