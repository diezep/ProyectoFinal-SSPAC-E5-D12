
module Ins_Mem(
input pcin,
output reg dataout
);
//Reg y wire
reg [31:0]insMem[31:0];

endmodule 