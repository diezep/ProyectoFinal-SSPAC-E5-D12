module modulo();



endmodule
